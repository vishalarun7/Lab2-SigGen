module counter #(
    parameter A_WIDTH = 8,
    parameter D_WIDTH = 8
)(
    //interface signals
    input logic clk, //clock
    input logic rst, //reset
    input logic en, //counter enable
    input logic [D_WIDTH-1:0] incr,
    output logic [A_WIDTH-1:0] count //count output 
);

always_ff @ (posedge clk)
    if (rst) count <= {A_WIDTH{1'b0}};
    else if (en) count <= count + incr;
endmodule
